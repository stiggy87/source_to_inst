// Verilog Test File 6

// Module #1

module 1st_module(port_1, port_2, port_3, port_4);
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
	
endmodule

// Module #2

module 2nd_module(port_1, port_2, port_3, port_4);
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
	
endmodule