// Verilog Test File 1

module test_1(port_1, port_2, port_3, port_4);
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
	
endmodule