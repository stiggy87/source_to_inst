// Verilog Test File 2

module test_2(
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
);

endmodule