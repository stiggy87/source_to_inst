// Verilog Test File 3

module test_3(
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
);

parameter WIDTH=6;
parameter HEIGHT=7;

endmodule