// Verilog Test File 5

module test_5
(
	input port_1,
	input port_2,
	inout port_3,
	output [1:0] port_4
);

endmodule