// Verilog Test File 4

module test_4(port_1, port_2, port_3, port_4);
	input port_1;
	input port_2;
	inout port_3;
	output [1:0] port_4;
	
	parameter WIDTH=6;
	parameter HEIGHT=7;
	
endmodule