entity test_1 is
	port (
		port_1 : in std_logic;
		port_2 : in std_logic;
		port_3 : inout std_logic;
		port_4 : out std_logic_vector (7 downto 0)
	);
end test_1;

